--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:56:40 04/08/2024
-- Design Name:   
-- Module Name:   /home/ise/Organosi/Ex1/mux8Tests.vhd
-- Project Name:  Ex1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: mux8
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY mux8Tests IS
END mux8Tests;
 
ARCHITECTURE behavior OF mux8Tests IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT mux8
    PORT(
         a1 : IN  std_logic_vector(31 downto 0);
         a2 : IN  std_logic_vector(31 downto 0);
         a3 : IN  std_logic_vector(31 downto 0);
         a4 : IN  std_logic_vector(31 downto 0);
         a5 : IN  std_logic_vector(31 downto 0);
         a6 : IN  std_logic_vector(31 downto 0);
         a7 : IN  std_logic_vector(31 downto 0);
         a8 : IN  std_logic_vector(31 downto 0);
         sel : IN  std_logic_vector(3 downto 0);
         b : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal a1 : std_logic_vector(31 downto 0) := (others => '0');
   signal a2 : std_logic_vector(31 downto 0) := (others => '0');
   signal a3 : std_logic_vector(31 downto 0) := (others => '0');
   signal a4 : std_logic_vector(31 downto 0) := (others => '0');
   signal a5 : std_logic_vector(31 downto 0) := (others => '0');
   signal a6 : std_logic_vector(31 downto 0) := (others => '0');
   signal a7 : std_logic_vector(31 downto 0) := (others => '0');
   signal a8 : std_logic_vector(31 downto 0) := (others => '0');
   signal sel : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal b : std_logic_vector(31 downto 0);
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: mux8 PORT MAP (
          a1 => a1,
          a2 => a2,
          a3 => a3,
          a4 => a4,
          a5 => a5,
          a6 => a6,
          a7 => a7,
          a8 => a8,
          sel => sel,
          b => b
        );

   -- Stimulus process
   stim_proc: process
   begin		
      wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "0000";
		wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "0001";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "0010";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "0011";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "0100";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "0101";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "0110";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "0111";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "1000";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "1001";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "1010";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "1011";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "1100";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "1101";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "1110";
		  wait for 10 ns;	
			a1 <= "00000000000000000000000000000000"; -- 0
			a2 <= "00000000000000000000000000000001"; -- 1
			a3 <= "00000000000000000000000000000010"; -- 2
			a4 <= "00000000000000000000000000000011"; -- 3
			a5 <= "00000000000000000000000000000100"; -- 4
			a6 <= "00000000000000000000000000000101"; -- 5
			a7 <= "00000000000000000000000000000110"; -- 6
			a8 <= "00000000000000000000000000000111"; -- 7
        sel <= "1111";
      -- insert stimulus here 

      wait;
   end process;

END;
